module tf_ROM 
    #(parameter addr_rom_width = 6,
                 data_width = 42,
                 depth_rom = 108)
    (
    input clk,
    input [addr_rom_width-1:0] A,
    input IREN,
    output reg [data_width-1:0] Q);
    
    always@(posedge clk)
    begin
    if(IREN == 1'b1) begin
    case(A)
    9'd0: Q <= 42'b011011111001111010100011101000111111001011;
    9'd1: Q <= 42'b001101110101101010101110100010100110010011;
    9'd2: Q <= 42'b101001100100110101100110100010001001010001;
    9'd3: Q <= 42'b100110000100000000101101001001011011100100;
    9'd4: Q <= 42'b001100011110110111111101101100100111110001;
    9'd5: Q <= 42'b001001000011110111010010110000110000010011;
    9'd6: Q <= 42'b100011100000001001011100000010010000010110;
    9'd7: Q <= 42'b101100010001100010100100111110110000011001;
    9'd8: Q <= 42'b010011110111101011000100110000101110010011;
    9'd9: Q <= 42'b001100000100110101100110000010001110000000;
    9'd10: Q <= 42'b100100011011100100111001111110101101101111;
    9'd11: Q <= 42'b011111001000010111100001001010101011010011;
    9'd12: Q <= 42'b100100000101100101101100010000001110111011;
    9'd13: Q <= 42'b010010111011101011011100111010111101110101;
    9'd14: Q <= 42'b010010110001011001000100001101111101100010;
    9'd15: Q <= 42'b100011110000101001000110001010110100101011;
    9'd16: Q <= 42'b101011110110111001010100100100011001100011;
    9'd17: Q <= 42'b101011011010001000110000000110001111000010;
    9'd18: Q <= 42'b101111011101010111001000111110001000100000;
    9'd19: Q <= 42'b101001100111100110010111000001110100010011;
    9'd20: Q <= 42'b011101111111100001010100011100010000100110;
    9'd21: Q <= 42'b001001011000010001001110110000100001110110;
    9'd22: Q <= 42'b000001100001100100100001100010111111111110;
    9'd23: Q <= 42'b011100000101000100010010010001110011001010;
    9'd24: Q <= 42'b100001000010000110011000011000000010100000;
    9'd25: Q <= 42'b000011111110010001111101110101110001001111;
    9'd26: Q <= 42'b000000000110110000101101100101110011100010;
    9'd27: Q <= 42'b000110011000001000110010100000101001010101;
    9'd28: Q <= 42'b100001010011100011001010100101101110110110;
    9'd29: Q <= 42'b000001011000100010010111101010101001101111;
    9'd30: Q <= 42'b010011100101000001011001010001001101001010;
    9'd31: Q <= 42'b100100101000010000010100111010100100010000;
    9'd32: Q <= 42'b001011001010110001101010000001101101010110;
    9'd33: Q <= 42'b000110000000010010110100000100111111011001;
    9'd34: Q <= 42'b100101100010110111000001110101111011000011;
    9'd35: Q <= 42'b010010011010100011001101010010001011011101;
    9'd36: Q <= 42'b010011100110111001111101100010011110000011;
    9'd37: Q <= 42'b001000011101101001001110011100001111111001;
    9'd38: Q <= 42'b101111011000010000111111111010000101001110;
    9'd39: Q <= 42'b101111100100000000011110000001110000100101;
    9'd40: Q <= 42'b101111111111100000000000100110111111100110;
    9'd41: Q <= 42'b001101001001001010010111100000000110000110;
    9'd42: Q <= 42'b100100111000100110110010111000000110111010;
    9'd43: Q <= 42'b001111110110010100001011011000111011000010;
    9'd44: Q <= 42'b001000011111100111001000010001001111101101;
    9'd45: Q <= 42'b001110001101001001100101110110010110001011;
    9'd46: Q <= 42'b101010011011110101101001111100000011110010;
    9'd47: Q <= 42'b010100101010110000010101001110110111100000;
    9'd48: Q <= 42'b000110011111110000100010000001110110010111;
    9'd49: Q <= 42'b011100010011110111111011000010010010100001;
    9'd50: Q <= 42'b010100010010110001010110010110011001010000;
    9'd51: Q <= 42'b001111110101011000100000000110111010011111;
    9'd52: Q <= 42'b011100111000101001100010010010010011010110;
    9'd53: Q <= 42'b000011111010101000011001001110011010100010;
    9'd54: Q <= 42'b011100100100011010010010001000101111001000;
    9'd55: Q <= 42'b010011111000000110111100011010001111000001;
    9'd56: Q <= 42'b100001001111011000011000011000101110111000;
    9'd57: Q <= 42'b101011110110000011100011010110011010111111;
    9'd58: Q <= 42'b000100100100000000001001000110010110000011;
    9'd59: Q <= 42'b101110011011010011011000001100110110110110;
    9'd60: Q <= 42'b101011010010100110100101101100111110001010;
    9'd61: Q <= 42'b100110011111000011010011011000111110010001;
    9'd62: Q <= 42'b100101111110111001100000110100000110100100;
    9'd63: Q <= 42'b010111100001101011101001111000000111011100;
    9'd64: Q <= 42'b011000011010100111110111101000100010000010;
    9'd65: Q <= 42'b000001111011011001010101011001010100011111;
    9'd66: Q <= 42'b011111000100000111001110011110010010111101;
    9'd67: Q <= 42'b011010101111011000001010010110100110100011;
    9'd68: Q <= 42'b000101011000100110001110101000100011001001;
    9'd69: Q <= 42'b100011010100101011000100100010011001111100;
    9'd70: Q <= 42'b100110101111110000110011101101100001101010;
    9'd71: Q <= 42'b100000011101111000010101110100101110101011;
    9'd72: Q <= 42'b010100110101000101101000011100101000000110;
    9'd73: Q <= 42'b100110101000100011110110110100010010010000;
    9'd74: Q <= 42'b100100010010010100010110010000100001011111;
    9'd75: Q <= 42'b011011101110101000110010000100110010110000;
    9'd76: Q <= 42'b001011110010000010010101110000000110010100;
    9'd77: Q <= 42'b000110010111100010011010110001001111100000;
    9'd78: Q <= 42'b101011100000000010001001010110100110111010;
    9'd79: Q <= 42'b010101000111110000000111011010110000010111;
    9'd80: Q <= 42'b100111001110000111000011011000111011000100;
    9'd81: Q <= 42'b011010010010100111101111111101101010111101;
    9'd82: Q <= 42'b001111100100010010110001010110111001001110;
    9'd83: Q <= 42'b100111011111110000001000001010111000010100;
    9'd84: Q <= 42'b001101110010110110110000001110101010011111;
    9'd85: Q <= 42'b000000000001110000000011000100000101010111;
    9'd86: Q <= 42'b001100010100100101110001101100010010111000;
    9'd87: Q <= 42'b000011010011010001001110111110100010001101;
    9'd88: Q <= 42'b001100110101010001011100101101010001011011;
    9'd89: Q <= 42'b001100001100000001011110100010101000000001;
    9'd90: Q <= 42'b100000100111001010001110101000001011001101;
    9'd91: Q <= 42'b011000001110110000010101111001111111111010;
    9'd92: Q <= 42'b001101110100000101010000011110101010100100;
    9'd93: Q <= 42'b000000110110001001100011110100001011001100;
    9'd94: Q <= 42'b000010111111111010011101001000100110010010;
    9'd95: Q <= 42'b011010011010111010100011000001101011011001;
    9'd96: Q <= 42'b100111010111000110001100101100000110100000;
    9'd97: Q <= 42'b001100100111010101001111100110001100110011;
    9'd98: Q <= 42'b000101000000101000110111111110111001001011;
    9'd99: Q <= 42'b101001010101111001111111100001101011011101;
    9'd100: Q <= 42'b000111111001010100011000110110101100111111;
    9'd101: Q <= 42'b100010011101000010111101011010000001111010;
    9'd102: Q <= 42'b010010010101010010010011100101111001101000;
    9'd103: Q <= 42'b011110101001100100000001001100110000001111;
    9'd104: Q <= 42'b100111000011001010001100111010101001111000;
    9'd105: Q <= 42'b101011000000010011110111101100101010011101;
    9'd106: Q <= 42'b101100011110010101111111111000100011010100;
    9'd107: Q <= 42'b101111111010010000100100000010101000000010;
    endcase end         
    end
endmodule